package ahb;

 `include "driver.sv"
 `include "generator.sv"
 `include "monitor.sv"
 `include "scoreboard.sv"

endpackage